wire clk;
pll u_pll(.clkin(clk_sys), .clkout0(clk));